module ImmGen (
    input logic [24:0] ImmInput,
    input logic [2:0] ImmSrc,

    output logic [31:0] ImmExt
);
    
endmodule